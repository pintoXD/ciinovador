module top;
   import uvm_pkg::*;
   import test_pkg::*;

   initial begin
      run_test("test");
   end
endmodule

