`include "uvm_macros.svh"
`include "bvm_macros.svh" // macros created by Brazil-IP / UFCG

package test_pkg;

  import uvm_pkg::*;

  `include "trans.svh"
  `include "source.svh"
  `include "refmod.svh"
  `include "sink.svh"
  `include "drain.svh"
  `include "env.svh"
  `include "test.svh"

endpackage
  
