class a_tr extends uvm_sequence_item;

  int a;

endclass

