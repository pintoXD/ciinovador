`include "uvm_macros.svh"
`include "bvm_macros.svh" // macros created by Brazil-IP / UFCG

package test_pkg;

  import uvm_pkg::*;

  `include "trans.svh"
  `include "source.svh"
  `include "sink.svh"
  `include "env.svh"
  `include "test.svh"

endpackage
  
