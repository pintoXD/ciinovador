module custom_ula(
    input logic [7:0] SrcA, SrcB,
    input logic [2:0] ULAControl,
    output logic [7:0] ULAResult,
    output logic FlagZ
);





endmodule custom_ula