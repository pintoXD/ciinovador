module notgate (a,b);
  input logic a;
  output logic b;
  
  assign b=!a;

endmodule